module test(
  input         clock,
  input         reset,
  input         io_valid,
  input  [63:0] io_bits_data,
  input  [63:0] io_bits_addr
);
endmodule
